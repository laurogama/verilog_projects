module somador ( input [3:0] a, b,

				output [4:0] c);
				
assign c = a + b;

endmodule
	